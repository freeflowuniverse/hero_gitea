module sub1

pub fn new2()! string{
	return "SSS2"
}