module vproto

import sub1

pub fn new()! string{
	println(sub1.new2()!)
	return "SSS"
}

